`timescale 1ns/1ns
module MUXnandTB();
logic aa,bb,cc,dd,s0,s1;
wire ww;
MUXnand CUT(aa,bb,cc,dd,s0,s1,ww);
initial begin
#20 aa=1;bb=0;cc=1;dd=0;
#50 s0=0;s1=0;
#50 s0=1;
#50 s1=0;
#50 s1=1;
#50 s0=1;
#50 s1=0;
#50 s0=0;
#50 s0=1;
#50 s1=1;
#50 s0=0;
#50 s1=0;
#50 aa=1;bb=0;cc=0;dd=1;
#50 s0=0;s1=0;
#50 s0=1;
#50 s1=0;
#50 s1=1;
#50 s0=1;
#50 s1=0;
#50 s0=0;
#50 s0=1;
#50 s1=1;
#50 s0=0;
#50 s1=0;
#50 $stop;
end
endmodule
