`timescale 1ns/1ns
module Bshifter16(input [15:0]A,[3:0]N,output [15:0]SHO);
MUX16to1 G1({A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15]},N,SHO[15]);
MUX16to1 G2({A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14]},N,SHO[14]);
MUX16to1 G3({A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13]},N,SHO[13]);
MUX16to1 G4({A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12]},N,SHO[12]);
MUX16to1 G5({A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11]},N,SHO[11]);
MUX16to1 G6({A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10]},N,SHO[10]);
MUX16to1 G7({A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9]},N,SHO[9]);
MUX16to1 G8({A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8]},N,SHO[8]);
MUX16to1 G9({A[6],A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7]},N,SHO[7]);
MUX16to1 G10({A[5],A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6]},N,SHO[6]);
MUX16to1 G11({A[4],A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5]},N,SHO[5]);
MUX16to1 G12({A[3],A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4]},N,SHO[4]);
MUX16to1 G13({A[2],A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3]},N,SHO[3]);
MUX16to1 G14({A[1],A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2]},N,SHO[2]);
MUX16to1 G15({A[0],A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1]},N,SHO[1]);
MUX16to1 G16({A[15],A[14],A[13],A[12],A[11],A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]},N,SHO[0]);
endmodule
